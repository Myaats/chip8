module cpu(input wire clk,
           input wire timer_cpu_tick,
           input wire timer_60hz_tick);
    
endmodule
