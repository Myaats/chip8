module cpu(input wire clk);

endmodule